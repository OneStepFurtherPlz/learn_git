module garb (  /*AUTOARG*/ );

  //=============================================================================
  //  parameter declare
  //=============================================================================


  //=============================================================================
  //  interface declare
  //=============================================================================
  /*AUTOTIEOFF*/
  input clk;    // Clock
  input rst_n;  // Asynchronous reset active low

  output [5:0] unused;


  input [4:0] dontcare;
  

  //=============================================================================
  //  wire/reg declaration
  //=============================================================================
  /*AUTOINPUT*/
  /*AUTOWIRE*/
  /*AUTOREG*/


endmodule
// Local Variables:
// verilog-auto-inst-param-value:t
// indent-tabs-mode:nil
// tab-width:2
// verilog-library-directories:(".")
// verilog-library-extensions:(".v")
// End:
