module test (  /*AUTOARG*/ );

  //=============================================================================
  //  parameter declare
  //=============================================================================


  //=============================================================================
  //  interface declare
  //=============================================================================
  /*AUTOTIEOFF*/
  input clk;    // Clock
  input rst_n;  // Asynchronous reset active low

  input [3:0] din;
  output [6 - 1: 0] dout;


  //=============================================================================
  //  wire/reg declaration
  //=============================================================================
  /*AUTOINPUT*/
  /*AUTOWIRE*/
  /*AUTOREG*/

  




endmodule
// Local Variables:
// verilog-auto-inst-param-value:t
// indent-tabs-mode:nil
// tab-width:2
// verilog-library-directories:(".")
// verilog-library-extensions:(".v")
// End:
